// Copyright 2020 Altera Corporation.
//
// This software and the related documents are Altera copyrighted materials,
// and your use of them is governed by the express license under which they
// were provided to you ("License"). Unless the License provides otherwise,
// you may not use, modify, copy, publish, distribute, disclose or transmit
// this software or the related documents without Altera's prior written
// permission.
//
// This software and the related documents are provided as is, with no express
// or implied warranties, other than those that are expressly stated in the
// License.

`resetall
`undefineall
`default_nettype none
`timescale 1ns/1ps

module dla_top_wrapper_AGX7_Generic_AGX7 #(
  // no input parameters needed
  //begining of autogenerated params
  localparam string DEVICE = "AGX7",
  localparam int C_CSR_AXI_ADDR_WIDTH = 11,
  localparam int C_CSR_AXI_DATA_WIDTH = 32,
  localparam int C_DDR_AXI_ADDR_WIDTH = 32,
  localparam int C_DDR_AXI_BURST_WIDTH = 4,
  localparam int C_DDR_AXI_DATA_WIDTH = 512,
  localparam int C_DDR_AXI_THREAD_ID_WIDTH = 2,
  localparam int CONFIG_DATA_BYTES = 4,
  localparam int CONFIG_READER_DATA_BYTES = 8,
  localparam int FILTER_READER_DATA_BYTES = 64,
  localparam int FEATURE_READER_DATA_BYTES = 32,
  localparam int FEATURE_WRITER_DATA_BYTES = 32,
  localparam int CONFIG_NUM_MODULES = 12,
  localparam int MODULE_ID_WIDTH = 8,
  localparam int CONFIG_CHANNEL_WIDTH = 32,
  localparam int CONFIG_CACHE_DEPTH = 256,
  localparam int CONFIG_NETWORK_QUANTIZE_DEPTHS [255:0] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,512,64,32},
  localparam bit CONFIG_NETWORK_CROSS_CLOCK [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,1},
  localparam bit CONFIG_NETWORK_CROSS_CLOCK_AXI [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
  localparam int CONFIG_NETWORK_FIFO_MIN_DEPTH [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256},
  localparam int CONFIG_NETWORK_NUM_PIPELINE_STAGES [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1},
  localparam int CONFIG_ID_PADDING = 0,
  localparam int CONFIG_ID_FILTER_READER = 1,
  localparam int CONFIG_ID_INPUT_FEEDER_MUX = 2,
  localparam int CONFIG_ID_INPUT_FEEDER_WRITER = 3,
  localparam int CONFIG_ID_INPUT_FEEDER_IN = 4,
  localparam int CONFIG_ID_INPUT_FEEDER_READER = 5,
  localparam int CONFIG_ID_INPUT_FEEDER_OUT = 6,
  localparam int CONFIG_ID_FEATURE_WRITER = 7,
  localparam int CONFIG_ID_FEATURE_READER = 8,
  localparam int CONFIG_ID_XBAR = 9,
  localparam int CONFIG_ID_ACTIVATION = 10,
  localparam int CONFIG_ID_POOL = 11,
  localparam int CONFIG_ID_SOFTMAX = 12,
  localparam bit ENABLE_DEBUG = 1,
  localparam bit ENABLE_INPUT_STREAMING = 0,
  localparam int AXI_ISTREAM_DATA_WIDTH = 128,
  localparam int AXI_ISTREAM_FIFO_DEPTH = 32,
  localparam bit ENABLE_ON_CHIP_PARAMETERS = 0,
  localparam bit ENABLE_MIXED_PRECISION = 0,
  localparam int KVEC_OVER_CVEC = 2,
  localparam int SB_ADDR_WIDTH = 16,
  localparam int STREAM_BUFFER_DEPTH = 63488,
  localparam bit[927:0] PE_ARRAY_PARAM_BITS = 928'h000000010000002000000001000000010000000900000009000000050000000f000000050000000f00000010000000030000000200000001000000010000000000000001000000000000000500000001000000020000000a00000004000000100000000000000001000000000000000100000003,
  localparam int PE_ARRAY_EXIT_FIFO_DEPTH = 1024,
  localparam int SCRATCHPAD_FILTER_DEPTH = 512,
  localparam int SCRATCHPAD_BIAS_SCALE_DEPTH = 512,
  localparam int SCRATCHPAD_NUM_FILTER_PORTS = 2,
  localparam int SCRATCHPAD_NUM_BIAS_SCALE_PORTS = 16,
  localparam int SCRATCHPAD_MEGABLOCK_WIDTH = 149,
  localparam int SCRATCHPAD_NUM_FILTER_BLOCKS_PER_MEGABLOCK = 1,
  localparam int SCRATCHPAD_NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK = 8,
  localparam int MAX_XBAR_INPUT_INTERFACES = 5,
  localparam int MAX_XBAR_OUTPUT_INTERFACES = 5,
  localparam int AUX_XBAR_INPUT_COUNTER_WIDTH = 24,
  localparam int AUX_XBAR_OUTPUT_COUNTER_WIDTH = 24,
  localparam bit ENABLE_ACTIVATION = 1,
  localparam bit ENABLE_DEPTHWISE = 0,
  localparam int XBAR_ID_DEPTHWISE = -1,
  localparam int CONFIG_ID_DEPTHWISE = -1,
  localparam bit ENABLE_DEPTHWISE_FILTER_BIAS = 0,
  localparam int XBAR_ID_DEPTHWISE_FILTER_BIAS = -1,
  localparam int CONFIG_ID_DEPTHWISE_FILTER_BIAS = -1,
  localparam bit ENABLE_POOL = 1,
  localparam bit ENABLE_SOFTMAX = 1,
  localparam int CONFIG_ID_OUTPUT_STREAMER = -1,
  localparam int CONFIG_ID_OUTPUT_STREAMER_FLUSH = -1,
  localparam int CONFIG_ID_WRITER_STREAMER_SEL = -1,
  localparam int CONFIG_ID_LAYOUT_TRANSFORM = -1,
  localparam int XBAR_ID_SOFTMAX = 3,
  localparam int XBAR_ID_POOL = 2,
  localparam int XBAR_ID_ACTIVATION = 1,
  localparam int XBAR_ID_XBAR_OUT_PORT = 0,
  localparam int XBAR_ID_PE_ARRAY = 0,
  localparam int NUMBER_OF_KERNELS = 3,
  localparam int AUX_MODULE_SELECT_ID_WIDTH = 4,
  localparam bit XBAR_KERNEL_BYPASS_FEATURE_ENABLE = 0,
  localparam bit AUX_KERNEL_BYPASSABLE [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0},
  localparam int AUX_XBAR_MUX_OUTPUT_PIPELINE_STAGES [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0},
  localparam int AUX_XBAR_NONSTALLABLE_OUTPUT_PIPELINE_STAGES [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0},
  localparam int AUX_XBAR_OUTPUT_BP_FIFO_ENABLE [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0},
  localparam int AUX_XBAR_OUTPUT_BP_FIFO_DEPTH [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0},
  localparam int AUX_XBAR_OUTPUT_WIDTH = 256,
  localparam int AUX_OUTPUT_DATA_WIDTHS [16:0] = '{0:256,1:256,2:256,3:256,4:256,5:256,6:256,7:256,8:256,9:256,10:256,11:256,12:256,13:256,14:256,15:256,16:256,default : 0},
  localparam int AUX_INPUT_DATA_WIDTHS [16:0] = '{0:256,1:256,2:256,3:256,4:256,5:256,6:256,7:256,8:256,9:256,10:256,11:256,12:256,13:256,14:256,15:256,16:256,default : 0},
  localparam int AUX_MAX_DATABUS_WIDTH = 256,
  localparam int XBAR_KERNEL_CV_FEATURE_ENABLE = 1,
  localparam int AUX_KERNEL_CONNECTIVITY_VECTOR [16:0] [16:0] = '{0: '{0:1,1:1,2:1,3:1,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},1: '{0:1,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},2: '{0:1,1:1,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},3: '{0:1,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},4: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},5: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},6: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},7: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},8: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},9: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},10: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},11: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},12: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},13: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},14: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},15: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},16: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0}},
  localparam int ACTIVATION_K_VECTOR = 16,
  localparam bit ACTIVATION_ENABLE_DSP_MULT = 0,
  localparam bit ACTIVATION_ENABLE_DSP_CONV = 0,
  localparam int ACTIVATION_GROUP_DELAY = 1,
  localparam int ACTIVATION_TYPE = 28,
  localparam int ACTIVATION_PARAM_CACHE_DEPTH = 1024,
  localparam int POOL_K_VECTOR = 4,
  localparam int POOL_GROUP_DELAY = 1,
  localparam int POOL_TYPE = 0,
  localparam int POOL_CONFIG_ID_WIDTH = 1,
  localparam int POOL_MAX_WINDOW_HEIGHT = 13,
  localparam int POOL_MAX_WINDOW_WIDTH = 13,
  localparam int POOL_MAX_STRIDE_VERTICAL = 4,
  localparam int POOL_MAX_STRIDE_HORIZONTAL = 4,
  localparam int POOL_PIPELINE_REG_NUM = 1,
  localparam int DEPTHWISE_K_VECTOR = 0,
  localparam int DEPTHWISE_GROUP_DELAY = 1,
  localparam int DEPTHWISE_TYPE = 0,
  localparam int DEPTHWISE_CONFIG_ID_WIDTH = 1,
  localparam int DEPTHWISE_MAX_WINDOW_HEIGHT = 3,
  localparam int DEPTHWISE_MAX_WINDOW_WIDTH = 3,
  localparam int DEPTHWISE_MAX_STRIDE_VERTICAL = 4,
  localparam int DEPTHWISE_MAX_STRIDE_HORIZONTAL = 4,
  localparam int DEPTHWISE_PIPELINE_REG_NUM = 1,
  localparam int DEPTHWISE_MAX_DILATION_VERTICAL = 1,
  localparam int DEPTHWISE_MAX_DILATION_HORIZONTAL = 1,
  localparam int DEPTHWISE_VECTOR_FEATURE_WIDTH = 16,
  localparam int DEPTHWISE_VECTOR_FILTER_WIDTH = 16,
  localparam int DEPTHWISE_VECTOR_BIAS_WIDTH = 32,
  localparam int DEPTHWISE_VECTOR_DOT_SIZE = 10,
  localparam int SOFTMAX_K_VECTOR = 1,
  localparam int SOFTMAX_GROUP_DELAY = 1,
  localparam int SOFTMAX_CONFIG_ID_WIDTH = 8,
  localparam int SOFTMAX_MAX_NUM_CHANNELS = 1024,
  localparam int AUX_MAX_TILE_HEIGHT = 128,
  localparam int AUX_MAX_TILE_WIDTH = 128,
  localparam int AUX_MAX_TILE_CHANNELS = 16384,
  localparam bit LAYOUT_TRANSFORM_ENABLE_IN_BIAS_SCALE = 0,
  localparam int LAYOUT_TRANSFORM_ENABLE = 0,
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_CHANNELS = 3,
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_HEIGHT = 28,
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_WIDTH = 28,
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_DEPTH = 1,
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_WIDTH = 2,
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_HEIGHT = 2,
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_DEPTH = 1,
  localparam int LAYOUT_TRANSFORM_MAX_PAD_FRONT = 1,
  localparam int LAYOUT_TRANSFORM_MAX_PAD_LEFT = 2,
  localparam int LAYOUT_TRANSFORM_MAX_PAD_TOP = 2,
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_HEIGHT = 2,
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_WIDTH = 2,
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_DEPTH = 1,
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_WIDTH = 2,
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_HEIGHT = 2,
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_DEPTH = 1,
  localparam int LAYOUT_TRANSFORM_READER_BYTES = 16,
  localparam int LAYOUT_TRANSFORM_DO_U8_CONV = 0,
  localparam int ENABLE_OUTPUT_STREAMER = 0,
  localparam int AXI_OSTREAM_DATA_WIDTH = 128,
  localparam int AXI_OSTREAM_ID_WIDTH = 8,
  localparam int AXI_OSTREAM_DEST_WIDTH = 8,
  localparam int AXI_OSTREAM_FIFO_DEPTH = 512,
  localparam int DISABLE_DDR = 0,
  //end of autogenerated params
  localparam int AXI_BURST_LENGTH_WIDTH = 8,  //width of the axi burst length signal as per the axi4 spec
  localparam int AXI_BURST_SIZE_WIDTH = 3,    //width of the axi burst size signal as per the axi4 spec
  localparam int AXI_BURST_TYPE_WIDTH = 2     //width of the axi burst type signal as per the axi4 spec
) (
  //clocks and resets, all resets are not synchronized
  input  wire                                     ddr_clk,
  input  wire                                     dla_clk,
  input  wire                                     axi_clk,
  input  wire                                     irq_clk,
  input  wire                                     dla_resetn,     //active low reset that has NOT been synchronized to any clock

  //interrupt request, AXI4 stream master without data, runs on pcie clock
  output logic                                    o_interrupt_level,

  //CSR, AXI4 lite slave, runs on ddr clock
  input  wire                                     i_csr_arvalid,
  input  wire          [C_CSR_AXI_ADDR_WIDTH-1:0] i_csr_araddr,
  output logic                                    o_csr_arready,
  output logic                                    o_csr_rvalid,
  output logic         [C_CSR_AXI_DATA_WIDTH-1:0] o_csr_rdata,
  input  wire                                     i_csr_rready,
  input  wire                                     i_csr_awvalid,
  input  wire          [C_CSR_AXI_ADDR_WIDTH-1:0] i_csr_awaddr,
  output logic                                    o_csr_awready,
  input  wire                                     i_csr_wvalid,
  input  wire          [C_CSR_AXI_DATA_WIDTH-1:0] i_csr_wdata,
  output logic                                    o_csr_wready,
  output logic                                    o_csr_bvalid,
  input  wire                                     i_csr_bready,

  //global memory, AXI4 master, runs on ddr clock
  output logic                                    o_ddr_arvalid,
  output logic         [C_DDR_AXI_ADDR_WIDTH-1:0] o_ddr_araddr,
  output logic       [AXI_BURST_LENGTH_WIDTH-1:0] o_ddr_arlen,
  output logic         [AXI_BURST_SIZE_WIDTH-1:0] o_ddr_arsize,
  output logic         [AXI_BURST_TYPE_WIDTH-1:0] o_ddr_arburst,
  output logic    [C_DDR_AXI_THREAD_ID_WIDTH-1:0] o_ddr_arid,
  input  wire                                     i_ddr_arready,
  input  wire                                     i_ddr_rvalid,
  input  wire          [C_DDR_AXI_DATA_WIDTH-1:0] i_ddr_rdata,
  input  wire     [C_DDR_AXI_THREAD_ID_WIDTH-1:0] i_ddr_rid,
  output logic                                    o_ddr_rready,
  output logic                                    o_ddr_awvalid,
  output logic         [C_DDR_AXI_ADDR_WIDTH-1:0] o_ddr_awaddr,
  output logic       [AXI_BURST_LENGTH_WIDTH-1:0] o_ddr_awlen,
  output logic         [AXI_BURST_SIZE_WIDTH-1:0] o_ddr_awsize,
  output logic         [AXI_BURST_TYPE_WIDTH-1:0] o_ddr_awburst,
  input  wire                                     i_ddr_awready,
  output logic                                    o_ddr_wvalid,
  output logic         [C_DDR_AXI_DATA_WIDTH-1:0] o_ddr_wdata,
  output logic     [(C_DDR_AXI_DATA_WIDTH/8)-1:0] o_ddr_wstrb,
  output logic                                    o_ddr_wlast,
  input  wire                                     i_ddr_wready,
  input  wire                                     i_ddr_bvalid,
  output logic                                    o_ddr_bready,

  // Input Streamer AXI-S interface signals
  input  wire                                     i_istream_axi_t_valid,
  output logic                                    o_istream_axi_t_ready,
  input  wire         [AXI_ISTREAM_DATA_WIDTH-1:0] i_istream_axi_t_data,

  // Output Streamer AXI-S interface signals
  output wire                                    o_ostream_axi_t_valid,
  input wire                                     i_ostream_axi_t_ready,
  output wire                                     o_ostream_axi_t_last,
  output logic   [AXI_OSTREAM_DATA_WIDTH-1:0]     o_ostream_axi_t_data,
  output logic   [(AXI_OSTREAM_DATA_WIDTH/8)-1:0] o_ostream_axi_t_strb
);

  dla_top #(
    .DEVICE                         (DEVICE),

    .CSR_ADDR_WIDTH                 (C_CSR_AXI_ADDR_WIDTH),
    .CSR_DATA_BYTES                 (C_CSR_AXI_DATA_WIDTH/8),
    .CONFIG_DATA_BYTES              (CONFIG_DATA_BYTES),
    .CONFIG_READER_DATA_BYTES       (CONFIG_READER_DATA_BYTES),
    .FILTER_READER_DATA_BYTES       (FILTER_READER_DATA_BYTES),
    .FEATURE_READER_DATA_BYTES      (FEATURE_READER_DATA_BYTES),
    .FEATURE_WRITER_DATA_BYTES      (FEATURE_WRITER_DATA_BYTES),
    .DDR_ADDR_WIDTH                 (C_DDR_AXI_ADDR_WIDTH),
    .DDR_DATA_BYTES                 (C_DDR_AXI_DATA_WIDTH/8),
    .DDR_BURST_WIDTH                (C_DDR_AXI_BURST_WIDTH),
    .DDR_READ_ID_WIDTH              (C_DDR_AXI_THREAD_ID_WIDTH),
    .ENABLE_ON_CHIP_PARAMETERS      (ENABLE_ON_CHIP_PARAMETERS),

    .KVEC_OVER_CVEC                 (KVEC_OVER_CVEC),
    .SB_ADDR_WIDTH                  (SB_ADDR_WIDTH),
    .STREAM_BUFFER_DEPTH            (STREAM_BUFFER_DEPTH),

    .PE_ARRAY_PARAM_BITS              (dla_pe_array_pkg::pe_array_arch_bits_t'(PE_ARRAY_PARAM_BITS)),
    .PE_ARRAY_EXIT_FIFO_DEPTH         (PE_ARRAY_EXIT_FIFO_DEPTH),

    .SCRATCHPAD_FILTER_DEPTH                       (SCRATCHPAD_FILTER_DEPTH),
    .SCRATCHPAD_BIAS_SCALE_DEPTH                   (SCRATCHPAD_BIAS_SCALE_DEPTH),
    .SCRATCHPAD_NUM_FILTER_PORTS                   (SCRATCHPAD_NUM_FILTER_PORTS),
    .SCRATCHPAD_NUM_BIAS_SCALE_PORTS               (SCRATCHPAD_NUM_BIAS_SCALE_PORTS),
    .SCRATCHPAD_MEGABLOCK_WIDTH                    (SCRATCHPAD_MEGABLOCK_WIDTH),
    .SCRATCHPAD_NUM_FILTER_BLOCKS_PER_MEGABLOCK    (SCRATCHPAD_NUM_FILTER_BLOCKS_PER_MEGABLOCK),
    .SCRATCHPAD_NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK(SCRATCHPAD_NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK),

    .CONFIG_NUM_MODULES             (CONFIG_NUM_MODULES),
    .MODULE_ID_WIDTH                (MODULE_ID_WIDTH),
    .CONFIG_CHANNEL_WIDTH           (CONFIG_CHANNEL_WIDTH),
    .CONFIG_CACHE_DEPTH             (CONFIG_CACHE_DEPTH),
    .CONFIG_ID_FILTER_READER        (CONFIG_ID_FILTER_READER),
    .CONFIG_ID_INPUT_FEEDER_MUX     (CONFIG_ID_INPUT_FEEDER_MUX),
    .CONFIG_ID_INPUT_FEEDER_WRITER  (CONFIG_ID_INPUT_FEEDER_WRITER),
    .CONFIG_ID_INPUT_FEEDER_IN      (CONFIG_ID_INPUT_FEEDER_IN),
    .CONFIG_ID_INPUT_FEEDER_READER  (CONFIG_ID_INPUT_FEEDER_READER),
    .CONFIG_ID_INPUT_FEEDER_OUT     (CONFIG_ID_INPUT_FEEDER_OUT),
    .CONFIG_ID_FEATURE_WRITER       (CONFIG_ID_FEATURE_WRITER),
    .CONFIG_ID_FEATURE_READER       (CONFIG_ID_FEATURE_READER),
    .CONFIG_ID_XBAR                 (CONFIG_ID_XBAR),
    .CONFIG_ID_OUTPUT_STREAMER      (CONFIG_ID_OUTPUT_STREAMER),
    .CONFIG_ID_OUTPUT_STREAMER_FLUSH(CONFIG_ID_OUTPUT_STREAMER_FLUSH),
    .CONFIG_ID_WRITER_STREAMER_SEL  (CONFIG_ID_WRITER_STREAMER_SEL),
    .CONFIG_ID_LAYOUT_TRANSFORM     (CONFIG_ID_LAYOUT_TRANSFORM),
    // AUX module config ID
    .CONFIG_ID_ACTIVATION           (CONFIG_ID_ACTIVATION),
    .CONFIG_ID_POOL                 (CONFIG_ID_POOL),
    .CONFIG_ID_DEPTHWISE            (CONFIG_ID_DEPTHWISE),
    .CONFIG_ID_DEPTHWISE_FILTER_BIAS(CONFIG_ID_DEPTHWISE_FILTER_BIAS),
    .CONFIG_ID_SOFTMAX              (CONFIG_ID_SOFTMAX),

    .CONFIG_NETWORK_QUANTIZE_DEPTHS (CONFIG_NETWORK_QUANTIZE_DEPTHS),
    .CONFIG_NETWORK_FIFO_MIN_DEPTH  (CONFIG_NETWORK_FIFO_MIN_DEPTH),
    .CONFIG_NETWORK_NUM_PIPELINE_STAGES (CONFIG_NETWORK_NUM_PIPELINE_STAGES),
    .CONFIG_NETWORK_CROSS_CLOCK     (CONFIG_NETWORK_CROSS_CLOCK),
    .CONFIG_NETWORK_CROSS_CLOCK_AXI (CONFIG_NETWORK_CROSS_CLOCK_AXI),

    //xbar
    .MAX_XBAR_INPUT_INTERFACES      (MAX_XBAR_INPUT_INTERFACES),
    .MAX_XBAR_OUTPUT_INTERFACES     (MAX_XBAR_OUTPUT_INTERFACES),
    .NUMBER_OF_KERNELS              (NUMBER_OF_KERNELS),
    .AUX_MODULE_SELECT_ID_WIDTH     (AUX_MODULE_SELECT_ID_WIDTH),
    .AUX_XBAR_INPUT_COUNTER_WIDTH   (AUX_XBAR_INPUT_COUNTER_WIDTH),
    .AUX_XBAR_OUTPUT_COUNTER_WIDTH  (AUX_XBAR_OUTPUT_COUNTER_WIDTH),
    .AUX_MAX_DATABUS_WIDTH          (AUX_MAX_DATABUS_WIDTH),
    .AUX_XBAR_OUTPUT_WIDTH          (AUX_XBAR_OUTPUT_WIDTH),
    .AUX_INPUT_DATA_WIDTHS          (AUX_INPUT_DATA_WIDTHS),
    .AUX_OUTPUT_DATA_WIDTHS         (AUX_OUTPUT_DATA_WIDTHS),
    .AUX_XBAR_MUX_OUTPUT_PIPELINE_STAGES(AUX_XBAR_MUX_OUTPUT_PIPELINE_STAGES),
    .AUX_XBAR_NONSTALLABLE_OUTPUT_PIPELINE_STAGES(AUX_XBAR_NONSTALLABLE_OUTPUT_PIPELINE_STAGES),
    .AUX_XBAR_OUTPUT_BP_FIFO_ENABLE (AUX_XBAR_OUTPUT_BP_FIFO_ENABLE),
    .AUX_XBAR_OUTPUT_BP_FIFO_DEPTH  (AUX_XBAR_OUTPUT_BP_FIFO_DEPTH),
    .XBAR_KERNEL_BYPASS_FEATURE_ENABLE (XBAR_KERNEL_BYPASS_FEATURE_ENABLE),
    .AUX_KERNEL_BYPASSABLE          (AUX_KERNEL_BYPASSABLE),
    .XBAR_KERNEL_CV_FEATURE_ENABLE  (XBAR_KERNEL_CV_FEATURE_ENABLE),
    .AUX_KERNEL_CONNECTIVITY_VECTOR (AUX_KERNEL_CONNECTIVITY_VECTOR),

    //xbar id
    .XBAR_ID_ACTIVATION             (XBAR_ID_ACTIVATION),
    .XBAR_ID_POOL                   (XBAR_ID_POOL),
    .XBAR_ID_DEPTHWISE              (XBAR_ID_DEPTHWISE),
    .XBAR_ID_SOFTMAX                (XBAR_ID_SOFTMAX),
    .XBAR_ID_PE_ARRAY               (XBAR_ID_PE_ARRAY),
    .XBAR_ID_XBAR_OUT_PORT          (XBAR_ID_XBAR_OUT_PORT),
    //aux module enable
    .ENABLE_ACTIVATION              (ENABLE_ACTIVATION),
    .ENABLE_POOL                    (ENABLE_POOL),
    .ENABLE_DEPTHWISE               (ENABLE_DEPTHWISE),
    .ENABLE_SOFTMAX                 (ENABLE_SOFTMAX),

    .ENABLE_INPUT_STREAMING         (ENABLE_INPUT_STREAMING),
    .AXI_ISTREAM_DATA_WIDTH         (AXI_ISTREAM_DATA_WIDTH),
    .AXI_ISTREAM_FIFO_DEPTH         (AXI_ISTREAM_FIFO_DEPTH),

    //debug module enable
    .ENABLE_DEBUG                   (ENABLE_DEBUG),

    // Output Streaming parameters
    .ENABLE_OUTPUT_STREAMER         (ENABLE_OUTPUT_STREAMER),
    .AXI_OSTREAM_DATA_WIDTH         (AXI_OSTREAM_DATA_WIDTH),
    .AXI_OSTREAM_ID_WIDTH           (AXI_OSTREAM_ID_WIDTH),
    .AXI_OSTREAM_DEST_WIDTH         (AXI_OSTREAM_DEST_WIDTH),
    .AXI_OSTREAM_FIFO_DEPTH         (AXI_OSTREAM_FIFO_DEPTH),

    // Mixed Precsion switch
    .ENABLE_MIXED_PRECISION         (ENABLE_MIXED_PRECISION),

    //Activation parameters
    .ACTIVATION_K_VECTOR            (ACTIVATION_K_VECTOR),
    .ACTIVATION_ENABLE_DSP_MULT     (ACTIVATION_ENABLE_DSP_MULT),
    .ACTIVATION_ENABLE_DSP_CONV     (ACTIVATION_ENABLE_DSP_CONV),
    .ACTIVATION_TYPE                (ACTIVATION_TYPE),
    .ACTIVATION_GROUP_DELAY         (ACTIVATION_GROUP_DELAY),
    .ACTIVATION_PARAM_CACHE_DEPTH   (ACTIVATION_PARAM_CACHE_DEPTH),

    //Pool parameters
    .POOL_K_VECTOR                  (POOL_K_VECTOR),
    .POOL_TYPE                      (POOL_TYPE),
    .POOL_GROUP_DELAY               (POOL_GROUP_DELAY),
    .POOL_CONFIG_ID_WIDTH           (POOL_CONFIG_ID_WIDTH),
    .POOL_MAX_WINDOW_HEIGHT         (POOL_MAX_WINDOW_HEIGHT),
    .POOL_MAX_WINDOW_WIDTH          (POOL_MAX_WINDOW_WIDTH),
    .POOL_MAX_STRIDE_VERTICAL       (POOL_MAX_STRIDE_VERTICAL),
    .POOL_MAX_STRIDE_HORIZONTAL     (POOL_MAX_STRIDE_HORIZONTAL),
    .POOL_PIPELINE_REG_NUM          (POOL_PIPELINE_REG_NUM),

    //Depthwise parameters
    .DEPTHWISE_K_VECTOR                  (DEPTHWISE_K_VECTOR),
    .DEPTHWISE_TYPE                      (DEPTHWISE_TYPE),
    .DEPTHWISE_GROUP_DELAY               (DEPTHWISE_GROUP_DELAY),
    .DEPTHWISE_CONFIG_ID_WIDTH           (DEPTHWISE_CONFIG_ID_WIDTH),
    .DEPTHWISE_MAX_WINDOW_HEIGHT         (DEPTHWISE_MAX_WINDOW_HEIGHT),
    .DEPTHWISE_MAX_WINDOW_WIDTH          (DEPTHWISE_MAX_WINDOW_WIDTH),
    .DEPTHWISE_MAX_STRIDE_VERTICAL       (DEPTHWISE_MAX_STRIDE_VERTICAL),
    .DEPTHWISE_MAX_STRIDE_HORIZONTAL     (DEPTHWISE_MAX_STRIDE_HORIZONTAL),
    .DEPTHWISE_PIPELINE_REG_NUM          (DEPTHWISE_PIPELINE_REG_NUM),
    .DEPTHWISE_MAX_DILATION_VERTICAL     (DEPTHWISE_MAX_DILATION_VERTICAL),
    .DEPTHWISE_MAX_DILATION_HORIZONTAL   (DEPTHWISE_MAX_DILATION_HORIZONTAL),

    // Depthwise vector parameters
    .DEPTHWISE_VECTOR_FEATURE_WIDTH      (DEPTHWISE_VECTOR_FEATURE_WIDTH),
    .DEPTHWISE_VECTOR_FILTER_WIDTH       (DEPTHWISE_VECTOR_FILTER_WIDTH),
    .DEPTHWISE_VECTOR_BIAS_WIDTH         (DEPTHWISE_VECTOR_BIAS_WIDTH),
    .DEPTHWISE_VECTOR_DOT_SIZE           (DEPTHWISE_VECTOR_DOT_SIZE),

    //Softmax parameters
    .SOFTMAX_K_VECTOR               (SOFTMAX_K_VECTOR),
    .SOFTMAX_GROUP_DELAY            (SOFTMAX_GROUP_DELAY),
    .SOFTMAX_CONFIG_ID_WIDTH        (SOFTMAX_CONFIG_ID_WIDTH),
    .SOFTMAX_MAX_NUM_CHANNELS       (SOFTMAX_MAX_NUM_CHANNELS),

    // Aux Parameters
    .AUX_MAX_TILE_HEIGHT            (AUX_MAX_TILE_HEIGHT),
    .AUX_MAX_TILE_WIDTH             (AUX_MAX_TILE_WIDTH),
    .AUX_MAX_TILE_CHANNELS             (AUX_MAX_TILE_CHANNELS),

    // Layout Transform
    .LAYOUT_TRANSFORM_ENABLE             (LAYOUT_TRANSFORM_ENABLE),
    .LAYOUT_TRANSFORM_ENABLE_IN_BIAS_SCALE   (LAYOUT_TRANSFORM_ENABLE_IN_BIAS_SCALE),
    .LAYOUT_TRANSFORM_MAX_FEATURE_CHANNELS   (LAYOUT_TRANSFORM_MAX_FEATURE_CHANNELS),
    .LAYOUT_TRANSFORM_MAX_FEATURE_HEIGHT     (LAYOUT_TRANSFORM_MAX_FEATURE_HEIGHT),
    .LAYOUT_TRANSFORM_MAX_FEATURE_WIDTH      (LAYOUT_TRANSFORM_MAX_FEATURE_WIDTH),
    .LAYOUT_TRANSFORM_MAX_FEATURE_DEPTH      (LAYOUT_TRANSFORM_MAX_FEATURE_DEPTH),
    .LAYOUT_TRANSFORM_MAX_STRIDE_WIDTH       (LAYOUT_TRANSFORM_MAX_STRIDE_WIDTH),
    .LAYOUT_TRANSFORM_MAX_STRIDE_HEIGHT      (LAYOUT_TRANSFORM_MAX_STRIDE_HEIGHT),
    .LAYOUT_TRANSFORM_MAX_STRIDE_DEPTH       (LAYOUT_TRANSFORM_MAX_STRIDE_DEPTH),
    .LAYOUT_TRANSFORM_MAX_PAD_FRONT          (LAYOUT_TRANSFORM_MAX_PAD_FRONT),
    .LAYOUT_TRANSFORM_MAX_PAD_LEFT           (LAYOUT_TRANSFORM_MAX_PAD_LEFT),
    .LAYOUT_TRANSFORM_MAX_PAD_TOP            (LAYOUT_TRANSFORM_MAX_PAD_TOP),
    .LAYOUT_TRANSFORM_MAX_FILTER_WIDTH       (LAYOUT_TRANSFORM_MAX_FILTER_WIDTH),
    .LAYOUT_TRANSFORM_MAX_FILTER_HEIGHT      (LAYOUT_TRANSFORM_MAX_FILTER_HEIGHT),
    .LAYOUT_TRANSFORM_MAX_FILTER_DEPTH       (LAYOUT_TRANSFORM_MAX_FILTER_DEPTH),
    .LAYOUT_TRANSFORM_MAX_DILATION_WIDTH     (LAYOUT_TRANSFORM_MAX_DILATION_WIDTH),
    .LAYOUT_TRANSFORM_MAX_DILATION_HEIGHT    (LAYOUT_TRANSFORM_MAX_DILATION_HEIGHT),
    .LAYOUT_TRANSFORM_MAX_DILATION_DEPTH     (LAYOUT_TRANSFORM_MAX_DILATION_DEPTH),
    .LAYOUT_TRANSFORM_READER_BYTES           (LAYOUT_TRANSFORM_READER_BYTES),
    .LAYOUT_TRANSFORM_DO_U8_CONV             (LAYOUT_TRANSFORM_DO_U8_CONV)
)
dla_top_inst
(
    .clk_ddr                        (ddr_clk),
    .clk_axi                        (axi_clk),
    .clk_dla                        (dla_clk),
    .clk_pcie                       (irq_clk),
    .i_resetn_async                 (dla_resetn),
    .o_interrupt_level              (o_interrupt_level),

    .i_csr_arvalid                  (i_csr_arvalid),
    .i_csr_araddr                   (i_csr_araddr),
    .o_csr_arready                  (o_csr_arready),
    .o_csr_rvalid                   (o_csr_rvalid),
    .o_csr_rdata                    (o_csr_rdata),
    .i_csr_rready                   (i_csr_rready),
    .i_csr_awvalid                  (i_csr_awvalid),
    .i_csr_awaddr                   (i_csr_awaddr),
    .o_csr_awready                  (o_csr_awready),
    .i_csr_wvalid                   (i_csr_wvalid),
    .i_csr_wdata                    (i_csr_wdata),
    .o_csr_wready                   (o_csr_wready),
    .o_csr_bvalid                   (o_csr_bvalid),
    .i_csr_bready                   (i_csr_bready),

    .o_ddr_arvalid                  (o_ddr_arvalid),
    .o_ddr_araddr                   (o_ddr_araddr),
    .o_ddr_arlen                    (o_ddr_arlen),
    .o_ddr_arsize                   (o_ddr_arsize),
    .o_ddr_arburst                  (o_ddr_arburst),
    .o_ddr_arid                     (o_ddr_arid),
    .i_ddr_arready                  (i_ddr_arready),
    .i_ddr_rvalid                   (i_ddr_rvalid),
    .i_ddr_rdata                    (i_ddr_rdata),
    .i_ddr_rid                      (i_ddr_rid),
    .o_ddr_rready                   (o_ddr_rready),
    .o_ddr_awvalid                  (o_ddr_awvalid),
    .o_ddr_awaddr                   (o_ddr_awaddr),
    .o_ddr_awlen                    (o_ddr_awlen),
    .o_ddr_awsize                   (o_ddr_awsize),
    .o_ddr_awburst                  (o_ddr_awburst),
    .i_ddr_awready                  (i_ddr_awready),
    .o_ddr_wvalid                   (o_ddr_wvalid),
    .o_ddr_wdata                    (o_ddr_wdata),
    .o_ddr_wstrb                    (o_ddr_wstrb),
    .o_ddr_wlast                    (o_ddr_wlast),
    .i_ddr_wready                   (i_ddr_wready),
    .i_ddr_bvalid                   (i_ddr_bvalid),
    .o_ddr_bready                   (o_ddr_bready),

    .i_istream_axi_t_valid          (i_istream_axi_t_valid),
    .o_istream_axi_t_ready          (o_istream_axi_t_ready),
    .i_istream_axi_t_data           (i_istream_axi_t_data),

    .o_ostream_axi_t_valid          (o_ostream_axi_t_valid),
    .i_ostream_axi_t_ready          (i_ostream_axi_t_ready),
    .o_ostream_axi_t_last           (o_ostream_axi_t_last),
    .o_ostream_axi_t_data           (o_ostream_axi_t_data),
    .o_ostream_axi_t_strb           (o_ostream_axi_t_strb)
);

endmodule
